module adder()
endmodule
